module top1 (inst_0_in2, inst_0_in1, inst_0_out1, inst_1_in3, inst_1_in2, inst_1_ctrl1, inst_1_out1, inst_2_in2, inst_2_in1, inst_2_out1, inst_3_in2, inst_3_in1, inst_3_out1, inst_4_in2, inst_4_in1, inst_4_out1, inst_5_in2, inst_5_ctrl1, inst_5_out1, inst_6_in2, inst_6_in1, inst_6_out1, inst_7_in2, inst_7_in1, inst_7_out1, inst_8_in2, inst_8_in1, inst_8_out1, inst_9_in2, inst_9_in1, inst_9_out1, inst_10_in2, inst_10_in1, inst_10_out1, inst_11_in2, inst_11_ctrl1, inst_11_out1, inst_12_in2, inst_12_in1, inst_12_out1, inst_13_in2, inst_13_in1, inst_13_out1, inst_14_in2, inst_14_in1, inst_14_out1, inst_15_in2, inst_15_in1, inst_15_out1, inst_16_in2, inst_16_in1, inst_16_out1, inst_17_in2, inst_17_in1, inst_17_out1, inst_18_in2, inst_18_in1, inst_18_out1, inst_19_in2, inst_19_in1, inst_19_out1, inst_20_in2, inst_20_in1, inst_20_out1, inst_21_in2, inst_21_in1, inst_21_out1, inst_22_in2, inst_22_in1, inst_22_out1, inst_23_in3, inst_23_in2, inst_23_ctrl1, inst_23_out1, inst_24_in1, inst_24_out1, inst_25_in2, inst_25_in1, inst_25_out1, inst_26_in2, inst_26_ctrl1, inst_26_out1, inst_27_in2, inst_27_in1, inst_27_out1, inst_28_in2, inst_28_in1, inst_28_out1, inst_29_in2, inst_29_in1, inst_29_out1, inst_30_in2, inst_30_in1, inst_30_out1, clk);

input [0:0] inst_0_in2;
wire [0:0] inst_0_in2_w;
reg [0:0] inst_0_in2_r;
input [0:0] inst_0_in1;
wire [0:0] inst_0_in1_w;
reg [0:0] inst_0_in1_r;
output [0:0] inst_0_out1;
wire [0:0] inst_0_out1_w;
reg [0:0] inst_0_out1_r;
input [0:0] inst_1_in3;
wire [0:0] inst_1_in3_w;
reg [0:0] inst_1_in3_r;
input [0:0] inst_1_in2;
wire [0:0] inst_1_in2_w;
reg [0:0] inst_1_in2_r;
input [0:0] inst_1_ctrl1;
wire [0:0] inst_1_ctrl1_w;
reg [0:0] inst_1_ctrl1_r;
output [0:0] inst_1_out1;
wire [0:0] inst_1_out1_w;
reg [0:0] inst_1_out1_r;
input [0:0] inst_2_in2;
wire [0:0] inst_2_in2_w;
reg [0:0] inst_2_in2_r;
input [0:0] inst_2_in1;
wire [0:0] inst_2_in1_w;
reg [0:0] inst_2_in1_r;
output [0:0] inst_2_out1;
wire [0:0] inst_2_out1_w;
reg [0:0] inst_2_out1_r;
input [31:0] inst_3_in2;
wire [31:0] inst_3_in2_w;
reg [31:0] inst_3_in2_r;
input [6:0] inst_3_in1;
wire [6:0] inst_3_in1_w;
reg [6:0] inst_3_in1_r;
output [31:0] inst_3_out1;
wire [31:0] inst_3_out1_w;
reg [31:0] inst_3_out1_r;
input [32:0] inst_4_in2;
wire [32:0] inst_4_in2_w;
reg [32:0] inst_4_in2_r;
input [31:0] inst_4_in1;
wire [31:0] inst_4_in1_w;
reg [31:0] inst_4_in1_r;
output [32:0] inst_4_out1;
wire [32:0] inst_4_out1_w;
reg [32:0] inst_4_out1_r;
input [31:0] inst_5_in2;
wire [31:0] inst_5_in2_w;
reg [31:0] inst_5_in2_r;
input [0:0] inst_5_ctrl1;
wire [0:0] inst_5_ctrl1_w;
reg [0:0] inst_5_ctrl1_r;
output [31:0] inst_5_out1;
wire [31:0] inst_5_out1_w;
reg [31:0] inst_5_out1_r;
input [31:0] inst_6_in2;
wire [31:0] inst_6_in2_w;
reg [31:0] inst_6_in2_r;
input [7:0] inst_6_in1;
wire [7:0] inst_6_in1_w;
reg [7:0] inst_6_in1_r;
output [0:0] inst_6_out1;
wire [0:0] inst_6_out1_w;
reg [0:0] inst_6_out1_r;
input [32:0] inst_7_in2;
wire [32:0] inst_7_in2_w;
reg [32:0] inst_7_in2_r;
input [32:0] inst_7_in1;
wire [32:0] inst_7_in1_w;
reg [32:0] inst_7_in1_r;
output [0:0] inst_7_out1;
wire [0:0] inst_7_out1_w;
reg [0:0] inst_7_out1_r;
input [31:0] inst_8_in2;
wire [31:0] inst_8_in2_w;
reg [31:0] inst_8_in2_r;
input [31:0] inst_8_in1;
wire [31:0] inst_8_in1_w;
reg [31:0] inst_8_in1_r;
output [0:0] inst_8_out1;
wire [0:0] inst_8_out1_w;
reg [0:0] inst_8_out1_r;
input [31:0] inst_9_in2;
wire [31:0] inst_9_in2_w;
reg [31:0] inst_9_in2_r;
input [1:0] inst_9_in1;
wire [1:0] inst_9_in1_w;
reg [1:0] inst_9_in1_r;
output [31:0] inst_9_out1;
wire [31:0] inst_9_out1_w;
reg [31:0] inst_9_out1_r;
input [6:0] inst_10_in2;
wire [6:0] inst_10_in2_w;
reg [6:0] inst_10_in2_r;
input [0:0] inst_10_in1;
wire [0:0] inst_10_in1_w;
reg [0:0] inst_10_in1_r;
output [6:0] inst_10_out1;
wire [6:0] inst_10_out1_w;
reg [6:0] inst_10_out1_r;
input [31:0] inst_11_in2;
wire [31:0] inst_11_in2_w;
reg [31:0] inst_11_in2_r;
input [0:0] inst_11_ctrl1;
wire [0:0] inst_11_ctrl1_w;
reg [0:0] inst_11_ctrl1_r;
output [31:0] inst_11_out1;
wire [31:0] inst_11_out1_w;
reg [31:0] inst_11_out1_r;
input [0:0] inst_12_in2;
wire [0:0] inst_12_in2_w;
reg [0:0] inst_12_in2_r;
input [0:0] inst_12_in1;
wire [0:0] inst_12_in1_w;
reg [0:0] inst_12_in1_r;
output [0:0] inst_12_out1;
wire [0:0] inst_12_out1_w;
reg [0:0] inst_12_out1_r;
input [31:0] inst_13_in2;
wire [31:0] inst_13_in2_w;
reg [31:0] inst_13_in2_r;
input [31:0] inst_13_in1;
wire [31:0] inst_13_in1_w;
reg [31:0] inst_13_in1_r;
output [0:0] inst_13_out1;
wire [0:0] inst_13_out1_w;
reg [0:0] inst_13_out1_r;
input [32:0] inst_14_in2;
wire [32:0] inst_14_in2_w;
reg [32:0] inst_14_in2_r;
input [1:0] inst_14_in1;
wire [1:0] inst_14_in1_w;
reg [1:0] inst_14_in1_r;
output [32:0] inst_14_out1;
wire [32:0] inst_14_out1_w;
reg [32:0] inst_14_out1_r;
input [31:0] inst_15_in2;
wire [31:0] inst_15_in2_w;
reg [31:0] inst_15_in2_r;
input [1:0] inst_15_in1;
wire [1:0] inst_15_in1_w;
reg [1:0] inst_15_in1_r;
output [31:0] inst_15_out1;
wire [31:0] inst_15_out1_w;
reg [31:0] inst_15_out1_r;
input [16:0] inst_16_in2;
wire [16:0] inst_16_in2_w;
reg [16:0] inst_16_in2_r;
input [0:0] inst_16_in1;
wire [0:0] inst_16_in1_w;
reg [0:0] inst_16_in1_r;
output [16:0] inst_16_out1;
wire [16:0] inst_16_out1_w;
reg [16:0] inst_16_out1_r;
input [12:0] inst_17_in2;
wire [12:0] inst_17_in2_w;
reg [12:0] inst_17_in2_r;
input [0:0] inst_17_in1;
wire [0:0] inst_17_in1_w;
reg [0:0] inst_17_in1_r;
output [12:0] inst_17_out1;
wire [12:0] inst_17_out1_w;
reg [12:0] inst_17_out1_r;
input [16:0] inst_18_in2;
wire [16:0] inst_18_in2_w;
reg [16:0] inst_18_in2_r;
input [31:0] inst_18_in1;
wire [31:0] inst_18_in1_w;
reg [31:0] inst_18_in1_r;
output [0:0] inst_18_out1;
wire [0:0] inst_18_out1_w;
reg [0:0] inst_18_out1_r;
input [31:0] inst_19_in2;
wire [31:0] inst_19_in2_w;
reg [31:0] inst_19_in2_r;
input [12:0] inst_19_in1;
wire [12:0] inst_19_in1_w;
reg [12:0] inst_19_in1_r;
output [31:0] inst_19_out1;
wire [31:0] inst_19_out1_w;
reg [31:0] inst_19_out1_r;
input [16:0] inst_20_in2;
wire [16:0] inst_20_in2_w;
reg [16:0] inst_20_in2_r;
input [32:0] inst_20_in1;
wire [32:0] inst_20_in1_w;
reg [32:0] inst_20_in1_r;
output [0:0] inst_20_out1;
wire [0:0] inst_20_out1_w;
reg [0:0] inst_20_out1_r;
input [15:0] inst_21_in2;
wire [15:0] inst_21_in2_w;
reg [15:0] inst_21_in2_r;
input [31:0] inst_21_in1;
wire [31:0] inst_21_in1_w;
reg [31:0] inst_21_in1_r;
output [0:0] inst_21_out1;
wire [0:0] inst_21_out1_w;
reg [0:0] inst_21_out1_r;
input [15:0] inst_22_in2;
wire [15:0] inst_22_in2_w;
reg [15:0] inst_22_in2_r;
input [0:0] inst_22_in1;
wire [0:0] inst_22_in1_w;
reg [0:0] inst_22_in1_r;
output [15:0] inst_22_out1;
wire [15:0] inst_22_out1_w;
reg [15:0] inst_22_out1_r;
input [31:0] inst_23_in3;
wire [31:0] inst_23_in3_w;
reg [31:0] inst_23_in3_r;
input [31:0] inst_23_in2;
wire [31:0] inst_23_in2_w;
reg [31:0] inst_23_in2_r;
input [0:0] inst_23_ctrl1;
wire [0:0] inst_23_ctrl1_w;
reg [0:0] inst_23_ctrl1_r;
output [31:0] inst_23_out1;
wire [31:0] inst_23_out1_w;
reg [31:0] inst_23_out1_r;
input [0:0] inst_24_in1;
wire [0:0] inst_24_in1_w;
reg [0:0] inst_24_in1_r;
output [0:0] inst_24_out1;
wire [0:0] inst_24_out1_w;
reg [0:0] inst_24_out1_r;
input [31:0] inst_25_in2;
wire [31:0] inst_25_in2_w;
reg [31:0] inst_25_in2_r;
input [31:0] inst_25_in1;
wire [31:0] inst_25_in1_w;
reg [31:0] inst_25_in1_r;
output [31:0] inst_25_out1;
wire [31:0] inst_25_out1_w;
reg [31:0] inst_25_out1_r;
input [31:0] inst_26_in2;
wire [31:0] inst_26_in2_w;
reg [31:0] inst_26_in2_r;
input [0:0] inst_26_ctrl1;
wire [0:0] inst_26_ctrl1_w;
reg [0:0] inst_26_ctrl1_r;
output [31:0] inst_26_out1;
wire [31:0] inst_26_out1_w;
reg [31:0] inst_26_out1_r;
input [31:0] inst_27_in2;
wire [31:0] inst_27_in2_w;
reg [31:0] inst_27_in2_r;
input [13:0] inst_27_in1;
wire [13:0] inst_27_in1_w;
reg [13:0] inst_27_in1_r;
output [0:0] inst_27_out1;
wire [0:0] inst_27_out1_w;
reg [0:0] inst_27_out1_r;
input [31:0] inst_28_in2;
wire [31:0] inst_28_in2_w;
reg [31:0] inst_28_in2_r;
input [1:0] inst_28_in1;
wire [1:0] inst_28_in1_w;
reg [1:0] inst_28_in1_r;
output [0:0] inst_28_out1;
wire [0:0] inst_28_out1_w;
reg [0:0] inst_28_out1_r;
input [31:0] inst_29_in2;
wire [31:0] inst_29_in2_w;
reg [31:0] inst_29_in2_r;
input [31:0] inst_29_in1;
wire [31:0] inst_29_in1_w;
reg [31:0] inst_29_in1_r;
output [31:0] inst_29_out1;
wire [31:0] inst_29_out1_w;
reg [31:0] inst_29_out1_r;
input [1:0] inst_30_in2;
wire [1:0] inst_30_in2_w;
reg [1:0] inst_30_in2_r;
input [31:0] inst_30_in1;
wire [31:0] inst_30_in1_w;
reg [31:0] inst_30_in1_r;
output [0:0] inst_30_out1;
wire [0:0] inst_30_out1_w;
reg [0:0] inst_30_out1_r;
input clk;

assign inst_0_in2_w = inst_0_in2_r;
assign inst_0_in1_w = inst_0_in1_r;
assign inst_0_out1 = inst_0_out1_r;
assign inst_1_in3_w = inst_1_in3_r;
assign inst_1_in2_w = inst_1_in2_r;
assign inst_1_ctrl1_w = inst_1_ctrl1_r;
assign inst_1_out1 = inst_1_out1_r;
assign inst_2_in2_w = inst_2_in2_r;
assign inst_2_in1_w = inst_2_in1_r;
assign inst_2_out1 = inst_2_out1_r;
assign inst_3_in2_w = inst_3_in2_r;
assign inst_3_in1_w = inst_3_in1_r;
assign inst_3_out1 = inst_3_out1_r;
assign inst_4_in2_w = inst_4_in2_r;
assign inst_4_in1_w = inst_4_in1_r;
assign inst_4_out1 = inst_4_out1_r;
assign inst_5_in2_w = inst_5_in2_r;
assign inst_5_ctrl1_w = inst_5_ctrl1_r;
assign inst_5_out1 = inst_5_out1_r;
assign inst_6_in2_w = inst_6_in2_r;
assign inst_6_in1_w = inst_6_in1_r;
assign inst_6_out1 = inst_6_out1_r;
assign inst_7_in2_w = inst_7_in2_r;
assign inst_7_in1_w = inst_7_in1_r;
assign inst_7_out1 = inst_7_out1_r;
assign inst_8_in2_w = inst_8_in2_r;
assign inst_8_in1_w = inst_8_in1_r;
assign inst_8_out1 = inst_8_out1_r;
assign inst_9_in2_w = inst_9_in2_r;
assign inst_9_in1_w = inst_9_in1_r;
assign inst_9_out1 = inst_9_out1_r;
assign inst_10_in2_w = inst_10_in2_r;
assign inst_10_in1_w = inst_10_in1_r;
assign inst_10_out1 = inst_10_out1_r;
assign inst_11_in2_w = inst_11_in2_r;
assign inst_11_ctrl1_w = inst_11_ctrl1_r;
assign inst_11_out1 = inst_11_out1_r;
assign inst_12_in2_w = inst_12_in2_r;
assign inst_12_in1_w = inst_12_in1_r;
assign inst_12_out1 = inst_12_out1_r;
assign inst_13_in2_w = inst_13_in2_r;
assign inst_13_in1_w = inst_13_in1_r;
assign inst_13_out1 = inst_13_out1_r;
assign inst_14_in2_w = inst_14_in2_r;
assign inst_14_in1_w = inst_14_in1_r;
assign inst_14_out1 = inst_14_out1_r;
assign inst_15_in2_w = inst_15_in2_r;
assign inst_15_in1_w = inst_15_in1_r;
assign inst_15_out1 = inst_15_out1_r;
assign inst_16_in2_w = inst_16_in2_r;
assign inst_16_in1_w = inst_16_in1_r;
assign inst_16_out1 = inst_16_out1_r;
assign inst_17_in2_w = inst_17_in2_r;
assign inst_17_in1_w = inst_17_in1_r;
assign inst_17_out1 = inst_17_out1_r;
assign inst_18_in2_w = inst_18_in2_r;
assign inst_18_in1_w = inst_18_in1_r;
assign inst_18_out1 = inst_18_out1_r;
assign inst_19_in2_w = inst_19_in2_r;
assign inst_19_in1_w = inst_19_in1_r;
assign inst_19_out1 = inst_19_out1_r;
assign inst_20_in2_w = inst_20_in2_r;
assign inst_20_in1_w = inst_20_in1_r;
assign inst_20_out1 = inst_20_out1_r;
assign inst_21_in2_w = inst_21_in2_r;
assign inst_21_in1_w = inst_21_in1_r;
assign inst_21_out1 = inst_21_out1_r;
assign inst_22_in2_w = inst_22_in2_r;
assign inst_22_in1_w = inst_22_in1_r;
assign inst_22_out1 = inst_22_out1_r;
assign inst_23_in3_w = inst_23_in3_r;
assign inst_23_in2_w = inst_23_in2_r;
assign inst_23_ctrl1_w = inst_23_ctrl1_r;
assign inst_23_out1 = inst_23_out1_r;
assign inst_24_in1_w = inst_24_in1_r;
assign inst_24_out1 = inst_24_out1_r;
assign inst_25_in2_w = inst_25_in2_r;
assign inst_25_in1_w = inst_25_in1_r;
assign inst_25_out1 = inst_25_out1_r;
assign inst_26_in2_w = inst_26_in2_r;
assign inst_26_ctrl1_w = inst_26_ctrl1_r;
assign inst_26_out1 = inst_26_out1_r;
assign inst_27_in2_w = inst_27_in2_r;
assign inst_27_in1_w = inst_27_in1_r;
assign inst_27_out1 = inst_27_out1_r;
assign inst_28_in2_w = inst_28_in2_r;
assign inst_28_in1_w = inst_28_in1_r;
assign inst_28_out1 = inst_28_out1_r;
assign inst_29_in2_w = inst_29_in2_r;
assign inst_29_in1_w = inst_29_in1_r;
assign inst_29_out1 = inst_29_out1_r;
assign inst_30_in2_w = inst_30_in2_r;
assign inst_30_in1_w = inst_30_in1_r;
assign inst_30_out1 = inst_30_out1_r;

mac_Xor_1Ux1U_1U_4 inst_0 (inst_0_in2_w, inst_0_in1_w, inst_0_out1_w);
mac_N_Muxb_1_2_4_4 inst_1 (inst_1_in3_w, inst_1_in2_w, inst_1_ctrl1_w, inst_1_out1_w);
mac_Or_1Ux1U_1U_4 inst_2 (inst_2_in2_w, inst_2_in1_w, inst_2_out1_w);
mac_Sub_32Sx7U_32S_4 inst_3 (inst_3_in2_w, inst_3_in1_w, inst_3_out1_w);
mac_Add_33Sx32U_33S_4 inst_4 (inst_4_in2_w, inst_4_in1_w, inst_4_out1_w);
mac_N_Mux_32_2_3_4 inst_5 (inst_5_in2_w, inst_5_ctrl1_w, inst_5_out1_w);
mac_GreaterThan_32Sx8S_1U_4 inst_6 (inst_6_in2_w, inst_6_in1_w, inst_6_out1_w);
mac_LessThan_33Sx33S_1U_4 inst_7 (inst_7_in2_w, inst_7_in1_w, inst_7_out1_w);
mac_LessThan_32Ux32U_1U_4 inst_8 (inst_8_in2_w, inst_8_in1_w, inst_8_out1_w);
mac_Add_32Sx2U_32S_4 inst_9 (inst_9_in2_w, inst_9_in1_w, inst_9_out1_w);
mac_Add_7Ux1U_7U_4 inst_10 (inst_10_in2_w, inst_10_in1_w, inst_10_out1_w);
mac_N_Mux_32_2_2_4 inst_11 (inst_11_in2_w, inst_11_ctrl1_w, inst_11_out1_w);
mac_And_1Ux1U_1U_4 inst_12 (inst_12_in2_w, inst_12_in1_w, inst_12_out1_w);
mac_Equal_32Ux32U_1U_4 inst_13 (inst_13_in2_w, inst_13_in1_w, inst_13_out1_w);
mac_Add_33Sx2U_33S_4 inst_14 (inst_14_in2_w, inst_14_in1_w, inst_14_out1_w);
mac_Add_32Ux2U_32U_4 inst_15 (inst_15_in2_w, inst_15_in1_w, inst_15_out1_w);
mac_Add_17Sx1U_17S_4 inst_16 (inst_16_in2_w, inst_16_in1_w, inst_16_out1_w);
mac_Add_13Sx1U_13S_4 inst_17 (inst_17_in2_w, inst_17_in1_w, inst_17_out1_w);
mac_LessThan_17Sx32S_1U_4 inst_18 (inst_18_in2_w, inst_18_in1_w, inst_18_out1_w);
mac_Sub_32Sx13U_32S_4 inst_19 (inst_19_in2_w, inst_19_in1_w, inst_19_out1_w);
mac_LessThan_17Sx33S_1U_4 inst_20 (inst_20_in2_w, inst_20_in1_w, inst_20_out1_w);
mac_LessThan_16Ux32U_1U_4 inst_21 (inst_21_in2_w, inst_21_in1_w, inst_21_out1_w);
mac_Add_16Ux1U_16U_4 inst_22 (inst_22_in2_w, inst_22_in1_w, inst_22_out1_w);
mac_N_MuxB_32_2_1_4 inst_23 (inst_23_in3_w, inst_23_in2_w, inst_23_ctrl1_w, inst_23_out1_w);
mac_Not_1U_1U_4 inst_24 (inst_24_in1_w, inst_24_out1_w);
mac_Add_32Ux32U_32U_4 inst_25 (inst_25_in2_w, inst_25_in1_w, inst_25_out1_w);
mac_N_Mux_32_2_0_4 inst_26 (inst_26_in2_w, inst_26_ctrl1_w, inst_26_out1_w);
mac_GreaterThan_32Sx14S_1U_4 inst_27 (inst_27_in2_w, inst_27_in1_w, inst_27_out1_w);
mac_GreaterThan_32Sx2S_1U_4 inst_28 (inst_28_in2_w, inst_28_in1_w, inst_28_out1_w);
mac_Mul_32Ux32U_32U_4 inst_29 (inst_29_in2_w, inst_29_in1_w, inst_29_out1_w);
mac_LessThan_2Sx32S_1U_4 inst_30 (inst_30_in2_w, inst_30_in1_w, inst_30_out1_w);

	always @ (posedge clk ) begin
		inst_0_in2_r <= inst_0_in2;
		inst_0_in1_r <= inst_0_in1;
		inst_0_out1_r <= inst_0_out1_w;
		inst_1_in3_r <= inst_1_in3;
		inst_1_in2_r <= inst_1_in2;
		inst_1_ctrl1_r <= inst_1_ctrl1;
		inst_1_out1_r <= inst_1_out1_w;
		inst_2_in2_r <= inst_2_in2;
		inst_2_in1_r <= inst_2_in1;
		inst_2_out1_r <= inst_2_out1_w;
		inst_3_in2_r <= inst_3_in2;
		inst_3_in1_r <= inst_3_in1;
		inst_3_out1_r <= inst_3_out1_w;
		inst_4_in2_r <= inst_4_in2;
		inst_4_in1_r <= inst_4_in1;
		inst_4_out1_r <= inst_4_out1_w;
		inst_5_in2_r <= inst_5_in2;
		inst_5_ctrl1_r <= inst_5_ctrl1;
		inst_5_out1_r <= inst_5_out1_w;
		inst_6_in2_r <= inst_6_in2;
		inst_6_in1_r <= inst_6_in1;
		inst_6_out1_r <= inst_6_out1_w;
		inst_7_in2_r <= inst_7_in2;
		inst_7_in1_r <= inst_7_in1;
		inst_7_out1_r <= inst_7_out1_w;
		inst_8_in2_r <= inst_8_in2;
		inst_8_in1_r <= inst_8_in1;
		inst_8_out1_r <= inst_8_out1_w;
		inst_9_in2_r <= inst_9_in2;
		inst_9_in1_r <= inst_9_in1;
		inst_9_out1_r <= inst_9_out1_w;
		inst_10_in2_r <= inst_10_in2;
		inst_10_in1_r <= inst_10_in1;
		inst_10_out1_r <= inst_10_out1_w;
		inst_11_in2_r <= inst_11_in2;
		inst_11_ctrl1_r <= inst_11_ctrl1;
		inst_11_out1_r <= inst_11_out1_w;
		inst_12_in2_r <= inst_12_in2;
		inst_12_in1_r <= inst_12_in1;
		inst_12_out1_r <= inst_12_out1_w;
		inst_13_in2_r <= inst_13_in2;
		inst_13_in1_r <= inst_13_in1;
		inst_13_out1_r <= inst_13_out1_w;
		inst_14_in2_r <= inst_14_in2;
		inst_14_in1_r <= inst_14_in1;
		inst_14_out1_r <= inst_14_out1_w;
		inst_15_in2_r <= inst_15_in2;
		inst_15_in1_r <= inst_15_in1;
		inst_15_out1_r <= inst_15_out1_w;
		inst_16_in2_r <= inst_16_in2;
		inst_16_in1_r <= inst_16_in1;
		inst_16_out1_r <= inst_16_out1_w;
		inst_17_in2_r <= inst_17_in2;
		inst_17_in1_r <= inst_17_in1;
		inst_17_out1_r <= inst_17_out1_w;
		inst_18_in2_r <= inst_18_in2;
		inst_18_in1_r <= inst_18_in1;
		inst_18_out1_r <= inst_18_out1_w;
		inst_19_in2_r <= inst_19_in2;
		inst_19_in1_r <= inst_19_in1;
		inst_19_out1_r <= inst_19_out1_w;
		inst_20_in2_r <= inst_20_in2;
		inst_20_in1_r <= inst_20_in1;
		inst_20_out1_r <= inst_20_out1_w;
		inst_21_in2_r <= inst_21_in2;
		inst_21_in1_r <= inst_21_in1;
		inst_21_out1_r <= inst_21_out1_w;
		inst_22_in2_r <= inst_22_in2;
		inst_22_in1_r <= inst_22_in1;
		inst_22_out1_r <= inst_22_out1_w;
		inst_23_in3_r <= inst_23_in3;
		inst_23_in2_r <= inst_23_in2;
		inst_23_ctrl1_r <= inst_23_ctrl1;
		inst_23_out1_r <= inst_23_out1_w;
		inst_24_in1_r <= inst_24_in1;
		inst_24_out1_r <= inst_24_out1_w;
		inst_25_in2_r <= inst_25_in2;
		inst_25_in1_r <= inst_25_in1;
		inst_25_out1_r <= inst_25_out1_w;
		inst_26_in2_r <= inst_26_in2;
		inst_26_ctrl1_r <= inst_26_ctrl1;
		inst_26_out1_r <= inst_26_out1_w;
		inst_27_in2_r <= inst_27_in2;
		inst_27_in1_r <= inst_27_in1;
		inst_27_out1_r <= inst_27_out1_w;
		inst_28_in2_r <= inst_28_in2;
		inst_28_in1_r <= inst_28_in1;
		inst_28_out1_r <= inst_28_out1_w;
		inst_29_in2_r <= inst_29_in2;
		inst_29_in1_r <= inst_29_in1;
		inst_29_out1_r <= inst_29_out1_w;
		inst_30_in2_r <= inst_30_in2;
		inst_30_in1_r <= inst_30_in1;
		inst_30_out1_r <= inst_30_out1_w;
	end
endmodule