module mux_64(out,sel,in0,in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16,in17,in18,in19,in20,in21,in22,in23,in24,in25,in26,in27,in28,in29,in30,in31,in32,in33,in34,in35,in36,in37,in38,in39,in40,in41,in42,in43,in44,in45,in46,in47,in48,in49,in50,in51,in52,in53,in54,in55,in56,in57,in58,in59,in60,in61,in62,in63);
output reg out;
input [5:0] sel;
input in0;
input in1;
input in2;
input in3;
input in4;
input in5;
input in6;
input in7;
input in8;
input in9;
input in10;
input in11;
input in12;
input in13;
input in14;
input in15;
input in16;
input in17;
input in18;
input in19;
input in20;
input in21;
input in22;
input in23;
input in24;
input in25;
input in26;
input in27;
input in28;
input in29;
input in30;
input in31;
input in32;
input in33;
input in34;
input in35;
input in36;
input in37;
input in38;
input in39;
input in40;
input in41;
input in42;
input in43;
input in44;
input in45;
input in46;
input in47;
input in48;
input in49;
input in50;
input in51;
input in52;
input in53;
input in54;
input in55;
input in56;
input in57;
input in58;
input in59;
input in60;
input in61;
input in62;
input in63;
always @(*) case (sel)
    0: out <= in0;
    1: out <= in1;
    2: out <= in2;
    3: out <= in3;
    4: out <= in4;
    5: out <= in5;
    6: out <= in6;
    7: out <= in7;
    8: out <= in8;
    9: out <= in9;
    10: out <= in10;
    11: out <= in11;
    12: out <= in12;
    13: out <= in13;
    14: out <= in14;
    15: out <= in15;
    16: out <= in16;
    17: out <= in17;
    18: out <= in18;
    19: out <= in19;
    20: out <= in20;
    21: out <= in21;
    22: out <= in22;
    23: out <= in23;
    24: out <= in24;
    25: out <= in25;
    26: out <= in26;
    27: out <= in27;
    28: out <= in28;
    29: out <= in29;
    30: out <= in30;
    31: out <= in31;
    32: out <= in32;
    33: out <= in33;
    34: out <= in34;
    35: out <= in35;
    36: out <= in36;
    37: out <= in37;
    38: out <= in38;
    39: out <= in39;
    40: out <= in40;
    41: out <= in41;
    42: out <= in42;
    43: out <= in43;
    44: out <= in44;
    45: out <= in45;
    46: out <= in46;
    47: out <= in47;
    48: out <= in48;
    49: out <= in49;
    50: out <= in50;
    51: out <= in51;
    52: out <= in52;
    53: out <= in53;
    54: out <= in54;
    55: out <= in55;
    56: out <= in56;
    57: out <= in57;
    58: out <= in58;
    59: out <= in59;
    60: out <= in60;
    61: out <= in61;
    62: out <= in62;
    63: out <= in63;
endcase
endmodule
