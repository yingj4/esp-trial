module top1 (inst_0_in3, inst_0_in2, inst_0_ctrl1, inst_0_out1, inst_1_in2, inst_1_in1, inst_1_out1, inst_2_in2, inst_2_in1, inst_2_out1, inst_3_in2, inst_3_in1, inst_3_out1, inst_4_in2, inst_4_in1, inst_4_out1, inst_5_in3, inst_5_in2, inst_5_ctrl1, inst_5_out1, inst_6_in2, inst_6_in1, inst_6_out1, inst_7_in2, inst_7_in1, inst_7_out1, inst_8_in2, inst_8_in1, inst_8_out1, clk);

input [31:0] inst_0_in3;
wire [31:0] inst_0_in3_w;
reg [31:0] inst_0_in3_r;
input [31:0] inst_0_in2;
wire [31:0] inst_0_in2_w;
reg [31:0] inst_0_in2_r;
input [0:0] inst_0_ctrl1;
wire [0:0] inst_0_ctrl1_w;
reg [0:0] inst_0_ctrl1_r;
output [31:0] inst_0_out1;
wire [31:0] inst_0_out1_w;
reg [31:0] inst_0_out1_r;
input [16:0] inst_1_in2;
wire [16:0] inst_1_in2_w;
reg [16:0] inst_1_in2_r;
input [1:0] inst_1_in1;
wire [1:0] inst_1_in1_w;
reg [1:0] inst_1_in1_r;
output [16:0] inst_1_out1;
wire [16:0] inst_1_out1_w;
reg [16:0] inst_1_out1_r;
input [13:0] inst_2_in2;
wire [13:0] inst_2_in2_w;
reg [13:0] inst_2_in2_r;
input [0:0] inst_2_in1;
wire [0:0] inst_2_in1_w;
reg [0:0] inst_2_in1_r;
output [13:0] inst_2_out1;
wire [13:0] inst_2_out1_w;
reg [13:0] inst_2_out1_r;
input [15:0] inst_3_in2;
wire [15:0] inst_3_in2_w;
reg [15:0] inst_3_in2_r;
input [1:0] inst_3_in1;
wire [1:0] inst_3_in1_w;
reg [1:0] inst_3_in1_r;
output [15:0] inst_3_out1;
wire [15:0] inst_3_out1_w;
reg [15:0] inst_3_out1_r;
input [12:0] inst_4_in2;
wire [12:0] inst_4_in2_w;
reg [12:0] inst_4_in2_r;
input [0:0] inst_4_in1;
wire [0:0] inst_4_in1_w;
reg [0:0] inst_4_in1_r;
output [12:0] inst_4_out1;
wire [12:0] inst_4_out1_w;
reg [12:0] inst_4_out1_r;
input [63:0] inst_5_in3;
wire [63:0] inst_5_in3_w;
reg [63:0] inst_5_in3_r;
input [63:0] inst_5_in2;
wire [63:0] inst_5_in2_w;
reg [63:0] inst_5_in2_r;
input [0:0] inst_5_ctrl1;
wire [0:0] inst_5_ctrl1_w;
reg [0:0] inst_5_ctrl1_r;
output [63:0] inst_5_out1;
wire [63:0] inst_5_out1_w;
reg [63:0] inst_5_out1_r;
input [31:0] inst_6_in2;
wire [31:0] inst_6_in2_w;
reg [31:0] inst_6_in2_r;
input [0:0] inst_6_in1;
wire [0:0] inst_6_in1_w;
reg [0:0] inst_6_in1_r;
output [31:0] inst_6_out1;
wire [31:0] inst_6_out1_w;
reg [31:0] inst_6_out1_r;
input [31:0] inst_7_in2;
wire [31:0] inst_7_in2_w;
reg [31:0] inst_7_in2_r;
input [0:0] inst_7_in1;
wire [0:0] inst_7_in1_w;
reg [0:0] inst_7_in1_r;
output [31:0] inst_7_out1;
wire [31:0] inst_7_out1_w;
reg [31:0] inst_7_out1_r;
input [31:0] inst_8_in2;
wire [31:0] inst_8_in2_w;
reg [31:0] inst_8_in2_r;
input [0:0] inst_8_in1;
wire [0:0] inst_8_in1_w;
reg [0:0] inst_8_in1_r;
output [31:0] inst_8_out1;
wire [31:0] inst_8_out1_w;
reg [31:0] inst_8_out1_r;
input clk;

assign inst_0_in3_w = inst_0_in3_r;
assign inst_0_in2_w = inst_0_in2_r;
assign inst_0_ctrl1_w = inst_0_ctrl1_r;
assign inst_0_out1 = inst_0_out1_r;
assign inst_1_in2_w = inst_1_in2_r;
assign inst_1_in1_w = inst_1_in1_r;
assign inst_1_out1 = inst_1_out1_r;
assign inst_2_in2_w = inst_2_in2_r;
assign inst_2_in1_w = inst_2_in1_r;
assign inst_2_out1 = inst_2_out1_r;
assign inst_3_in2_w = inst_3_in2_r;
assign inst_3_in1_w = inst_3_in1_r;
assign inst_3_out1 = inst_3_out1_r;
assign inst_4_in2_w = inst_4_in2_r;
assign inst_4_in1_w = inst_4_in1_r;
assign inst_4_out1 = inst_4_out1_r;
assign inst_5_in3_w = inst_5_in3_r;
assign inst_5_in2_w = inst_5_in2_r;
assign inst_5_ctrl1_w = inst_5_ctrl1_r;
assign inst_5_out1 = inst_5_out1_r;
assign inst_6_in2_w = inst_6_in2_r;
assign inst_6_in1_w = inst_6_in1_r;
assign inst_6_out1 = inst_6_out1_r;
assign inst_7_in2_w = inst_7_in2_r;
assign inst_7_in1_w = inst_7_in1_r;
assign inst_7_out1 = inst_7_out1_r;
assign inst_8_in2_w = inst_8_in2_r;
assign inst_8_in1_w = inst_8_in1_r;
assign inst_8_out1 = inst_8_out1_r;

mac_N_Mux_32_2_2_4 inst_0 (inst_0_in3_w, inst_0_in2_w, inst_0_ctrl1_w, inst_0_out1_w);
mac_Add_17Sx2U_17S_4 inst_1 (inst_1_in2_w, inst_1_in1_w, inst_1_out1_w);
mac_Add_14Sx1U_14S_4 inst_2 (inst_2_in2_w, inst_2_in1_w, inst_2_out1_w);
mac_Add_16Ux2U_16U_4 inst_3 (inst_3_in2_w, inst_3_in1_w, inst_3_out1_w);
mac_Add_13Ux1U_13U_4 inst_4 (inst_4_in2_w, inst_4_in1_w, inst_4_out1_w);
mac_N_MuxB_64_2_1_4 inst_5 (inst_5_in3_w, inst_5_in2_w, inst_5_ctrl1_w, inst_5_out1_w);
mac_Add_32Sx1U_32S_4 inst_6 (inst_6_in2_w, inst_6_in1_w, inst_6_out1_w);
mac_Or_32Sx1U_32S_4 inst_7 (inst_7_in2_w, inst_7_in1_w, inst_7_out1_w);
mac_Sub_32Sx1U_32S_4 inst_8 (inst_8_in2_w, inst_8_in1_w, inst_8_out1_w);

	always @ (posedge clk ) begin
		inst_0_in3_r <= inst_0_in3;
		inst_0_in2_r <= inst_0_in2;
		inst_0_ctrl1_r <= inst_0_ctrl1;
		inst_0_out1_r <= inst_0_out1_w;
		inst_1_in2_r <= inst_1_in2;
		inst_1_in1_r <= inst_1_in1;
		inst_1_out1_r <= inst_1_out1_w;
		inst_2_in2_r <= inst_2_in2;
		inst_2_in1_r <= inst_2_in1;
		inst_2_out1_r <= inst_2_out1_w;
		inst_3_in2_r <= inst_3_in2;
		inst_3_in1_r <= inst_3_in1;
		inst_3_out1_r <= inst_3_out1_w;
		inst_4_in2_r <= inst_4_in2;
		inst_4_in1_r <= inst_4_in1;
		inst_4_out1_r <= inst_4_out1_w;
		inst_5_in3_r <= inst_5_in3;
		inst_5_in2_r <= inst_5_in2;
		inst_5_ctrl1_r <= inst_5_ctrl1;
		inst_5_out1_r <= inst_5_out1_w;
		inst_6_in2_r <= inst_6_in2;
		inst_6_in1_r <= inst_6_in1;
		inst_6_out1_r <= inst_6_out1_w;
		inst_7_in2_r <= inst_7_in2;
		inst_7_in1_r <= inst_7_in1;
		inst_7_out1_r <= inst_7_out1_w;
		inst_8_in2_r <= inst_8_in2;
		inst_8_in1_r <= inst_8_in1;
		inst_8_out1_r <= inst_8_out1_w;
	end
endmodule