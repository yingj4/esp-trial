/*****************************************************************************
    Verilog RTL Description
    
    Configured at: 16:21:48 CDT (-0500), Sunday 28 March 2021
    Configured on: mojave.cs.illinois.edu
    Configured by: yingj4 (Ying Jing)
    
    Created by: Stratus DpOpt 2019.1.02 
*******************************************************************************/

module mac_LessThan_2Sx32S_1U_4 (
	in2,
	in1,
	out1
	); /* architecture "behavioural" */ 
input [1:0] in2;
input [31:0] in1;
output  out1;
wire  asc001;

assign asc001 = ($signed(in1)>$signed(in2));

assign out1 = asc001;
endmodule

/* CADENCE  urn3Qw0= : u9/ySgnWtBlWxVDRXgAb5+g= ** DO NOT EDIT THIS LINE ******/

